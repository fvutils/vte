/****************************************************************************
 * {{name}}_seq_item.svh
 * 
 ****************************************************************************/
{% set filename = "{{name}}_seq_item.svh" %} 

class {{name}}_seq_item `{{name}}_plist extends uvm_sequence_item;
	typedef {{name}}_seq_item `{{name}}_params this_t;
	`uvm_object_param_utils(this_t)
	
	const string report_id = "{{name}}_seq_item";
	
	// TODO: Declare fields here
	
	function new(string name="{{name}}_seq_item");
		super.new(name);
	endfunction

	// TODO: Declare do_print, do_compare, do_copy methods

	function void do_print(uvm_printer printer);
		if (printer.knobs.sprint == 0) begin
			$display(convert2string());
		end else begin
			printer.m_string = convert2string();
		end
	endfunction

	function bit do_compare(uvm_object rhs, uvm_comparer comparer);
		bit ret = 1;
		{{name}}_seq_item rhs_;
		
		if (!$cast(rhs_, rhs)) begin
			return 0;
		end
		
		ret &= super.do_compare(rhs, comparer);
		
		// TODO: implement comparison logic
	
		return ret;
	endfunction

	function void do_copy(uvm_object rhs);
		{{name}}_seq_item rhs_;
		
		if (!$cast(rhs_, rhs)) begin
			`uvm_error(report_id, "Cast failed in do_copy()");
			return;
		end
		
		super.do_copy(rhs);
		
		// TODO: copy item-specific fields
		
	endfunction
			
endclass



