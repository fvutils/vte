
{%set filename = "tests/{{name}}_tests_pkg.sv" %}

`include "uvm_macros.svh"
package {{name}}_tests_pkg;
	import uvm_pkg::*;
	import {{name}}_env_pkg::*;
	
	`include "{{name}}_test_base.svh"
	
endpackage
